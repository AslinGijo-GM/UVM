interface intf(input clk);
   
	logic clk;
   logic[3:0] A;
   logic[3:0] B;
  logic [5:0] Result;
   logic [2:0] sel;
  
  
   
  
endinterface 

interface intf(input logic clk,reset);
  
 // logic clk   ;
  logic d     ;
 // logic reset ;
  logic q     ;
  
endinterface
